//module sigma_tb;


//reg clk;
//reg reset_n;
//reg [31:0] A00, A01, A02;
//reg [31:0] A10, A11, A12;
//reg [31:0] A20, A21, A22;
//wire [31:0] sigma;
//wire valid;

//sigma#(
//	.PRECISION(32)
//) uut(
//	.clk(clk), .reset_n(reset_n),
//	.err(32'h3dcccccd),
//	.A00(A00), .A01(A01), .A02(A02),
//	.A10(A10), .A11(A11), .A12(A12),
//	.A20(A20), .A21(A21), .A22(A22),
//	.valid(valid),
//	.sigma(sigma)
//);

//initial begin
//    	clk = 0;
//    	forever #5 clk = ~clk;
//end

//initial begin
//    	reset_n   = 0;

//    	#25;
//    	reset_n = 1;

//    	@(posedge clk);
//        A00 <= 0;
//        A01 <= 32'h3f000000;
//        A02 <= 32'h3d4ccccd;
    
//        A10 <= 32'h3eaaaaaa;
//        A11 <= 0;
//        A12 <= 32'h3eaaaaaa;
    
//        A20 <= 32'h3d4ccccd;
//        A21 <= 32'h3f000000;
//        A22 <= 0;
//        #2000;

//    	$finish;
//end
//endmodule

module sigma_tb;

reg clk;
reg reset_n;
reg [31:0] A00, A01, A02;
reg [31:0] A10, A11, A12;
reg [31:0] A20, A21, A22;
wire [31:0] sigma;
wire valid;

integer cycle_count;
integer start_cycle, end_cycle;
real clk_period = 10.0; // 10ns = 100MHz

sigma#(
	.PRECISION(32)
) uut(
	.clk(clk), .reset_n(reset_n),
	.err(32'h3dcccccd),
	.A00(A00), .A01(A01), .A02(A02),
	.A10(A10), .A11(A11), .A12(A12),
	.A20(A20), .A21(A21), .A22(A22),
	.valid(valid),
	.sigma(sigma)
);

// Clock
initial begin
    	clk = 0;
    	forever #5 clk = ~clk; // 100MHz
end

// Stimulus
initial begin
    	reset_n = 0;
    	#25;
    	reset_n = 1;

    	@(posedge clk);
    	A00 <= 0;
    	A01 <= 32'h3f000000;
    	A02 <= 32'h3d4ccccd;

    	A10 <= 32'h3eaaaaaa;
    	A11 <= 0;
    	A12 <= 32'h3eaaaaaa;

    	A20 <= 32'h3d4ccccd;
    	A21 <= 32'h3f000000;
    	A22 <= 0;

    	start_cycle = cycle_count; // bắt đầu đếm
    	
    	wait(valid == 1'b1); // chờ đến khi output hợp lệ
    	end_cycle = cycle_count;

    	$display("\n===========================================");
    	$display("Sigma output = %h", sigma);
    	$display("Latency = %0d cycles", end_cycle - start_cycle);
    	$display("Latency = %.1f ns", (end_cycle - start_cycle) * clk_period);
    	$display("===========================================\n");

    	#50;
    	$finish;
end

// Cycle counter
always @(posedge clk or negedge reset_n) begin
	if (!reset_n)
		cycle_count <= 0;
	else
		cycle_count <= cycle_count + 1;
end

endmodule
