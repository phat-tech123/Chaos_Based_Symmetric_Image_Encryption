module Crypto_Engine_top();



endmodule
